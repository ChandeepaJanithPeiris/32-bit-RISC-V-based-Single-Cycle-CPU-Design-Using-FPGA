library verilog;
use verilog.vl_types.all;
entity program_counter_tb is
end program_counter_tb;
